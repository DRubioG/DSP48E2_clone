library ieee;
use ieee.std_logic_11